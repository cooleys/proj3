//-----------------------------------------------------------------------------
// Title         : MIPS Single-Cycle Control Unit
// Project       : ECE 313 - Computer Organization
//-----------------------------------------------------------------------------
// File          : control_single.v
// Author        : John Nestor  <nestorj@lafayette.edu>
// Organization  : Lafayette College
// 
// Created       : October 2002
// Last modified : 7 January 2005
//-----------------------------------------------------------------------------
// Description :
//   Control unit for the MIPS "Single Cycle" processor implementation described
//   Section 5.4 of "Computer Organization and Design, 3rd ed."
//   by David Patterson & John Hennessey, Morgan Kaufmann, 2004 (COD3e).  
//
//   It implements the function specified in Figure 5.18 on p. 308 of COD3e.
//
//-----------------------------------------------------------------------------

module control_single(opcode, RegDst, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, BranchNE, Jump, ALUOp);
    input [5:0] opcode;

	// Add Jump and BranchNE to the optputs
    output RegDst, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, BranchNE, Jump;
    output [1:0] ALUOp;
    reg    RegDst, ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch, BranchNE, Jump;
    reg    [1:0] ALUOp;

	// Add J, ADDI, and BNE to our instructions and codes
    parameter R_FORMAT = 6'd0;
    parameter LW = 6'd35;
    parameter SW = 6'd43;
    parameter BEQ = 6'd4;
	parameter BNE = 6'd5;
	parameter J = 6'd2;
	parameter ADDI = 6'd8;

    always @(opcode)
    begin
        case (opcode)
          R_FORMAT : 
          begin
              RegDst=1'b1;
			  ALUSrc=1'b0;
			  MemtoReg=1'b0; 
			  RegWrite=1'b1; 
			  MemRead=1'b0; 
              MemWrite=1'b0;
			  Branch=1'b0;
			  BranchNE = 1'b0;
			  Jump = 1'b0;
			  ALUOp = 2'b10;
          end
          
		  LW :
          begin
              RegDst=1'b0;
			  ALUSrc=1'b1; 
			  MemtoReg=1'b1;
			  RegWrite=1'b1;
			  MemRead=1'b1; 
              MemWrite=1'b0; 
			  Branch=1'b0; 
			  BranchNE = 1'b0;
			  Jump = 1'b0;
			  ALUOp = 2'b00;
          end
          
		  SW :
          begin
              RegDst=1'bx;
			  ALUSrc=1'b1;
			  MemtoReg=1'bx;
			  RegWrite=1'b0;
			  MemRead=1'b0; 
              MemWrite=1'b1;
			  Branch=1'b0;
			  BranchNE = 1'b0;
			  Jump = 1'b0;
			  ALUOp = 2'b00;
          end
          
		  BEQ :
          begin
              RegDst=1'bx;
			  ALUSrc=1'b0; 
			  MemtoReg=1'bx; 
			  RegWrite=1'b0; 
			  MemRead=1'b0; 
              MemWrite=1'b0; 
			  Branch=1'b1; 
			  BranchNE = 1'b0;
			  Jump = 1'b0;
			  ALUOp = 2'b01;
          end

		 BNE :
		 begin
		 	RegDst=1'bx;
			ALUSrc=1'b0; 
			MemtoReg=1'bx; 
			RegWrite=1'b0; 
			MemRead=1'b0; 
            MemWrite=1'b0; 
			Branch=1'b0; 
			BranchNE = 1'b1;
			Jump = 1'b0;
			ALUOp = 2'b01;
		  end

		  J :
		  begin
		 	RegDst=1'bx;
			ALUSrc=1'b0; 
			MemtoReg=1'bx; 
			RegWrite=1'bx; 
			MemRead=1'bx; 
            MemWrite=1'bx; 
			Branch=1'b1; 
			BranchNE = 1'b0;
			Jump = 1'b1;
			ALUOp = 2'b01;
		  	
		  end

		  ADDI :
		  begin
		 	RegDst=1'b1;
			ALUSrc=1'b0; 
			MemtoReg=1'b0; 
			RegWrite=1'b1; 
			MemRead=1'b0; 
            MemWrite=1'b0; 
			Branch=1'b0; 
			BranchNE = 1'b0;
			Jump = 1'b0;
			ALUOp = 2'b10;	
		  end

          default
          begin
              $display("control_single unimplemented opcode %d", opcode);
              RegDst=1'bx; ALUSrc=1'bx; MemtoReg=1'bx; RegWrite=1'bx; MemRead=1'bx; 
              MemWrite=1'bx; Branch=1'bx; ALUOp = 2'bxx;
          end

        endcase
    end
endmodule

